--reciprocal.vhd
-- Generated at Mon Aug 13 12:50:23 2018
--Andrew Miller 8/13/18
--reciprocal.vhd is a 32 bit reicprocal approximator

library IEEE;
use IEEE.std_logic_1164.all;

entity reciprocal is

  port(
       b : in std_logic_vector(31 downto 0);
       r : out std_logic_vector(31 downto 0)
       );
  
end entity reciprocal;

architecture default of reciprocal is

  
begin

  r <= "11000000000000000000000000000000" when b               = "00000000000000000000000000000000" else
       "01100000000000000000000000000000" when b(31 downto 1)  = "0000000000000000000000000000000" else
       "00110000000000000000000000000000" when b(31 downto 2)  = "000000000000000000000000000000" else
       "00011000000000000000000000000000" when b(31 downto 3)  = "00000000000000000000000000000" else
       "00001100000000000000000000000000" when b(31 downto 4)  = "0000000000000000000000000000" else
       "00000110000000000000000000000000" when b(31 downto 5)  = "000000000000000000000000000" else
       "00000011000000000000000000000000" when b(31 downto 6)  = "00000000000000000000000000" else
       "00000001100000000000000000000000" when b(31 downto 7)  = "0000000000000000000000000" else
       "00000000110000000000000000000000" when b(31 downto 8)  = "000000000000000000000000" else
       "00000000011000000000000000000000" when b(31 downto 9)  = "00000000000000000000000" else
       "00000000001100000000000000000000" when b(31 downto 10) = "0000000000000000000000" else
       "00000000000110000000000000000000" when b(31 downto 11) = "000000000000000000000" else
       "00000000000011000000000000000000" when b(31 downto 12) = "00000000000000000000" else
       "00000000000001100000000000000000" when b(31 downto 13) = "0000000000000000000" else
       "00000000000000110000000000000000" when b(31 downto 14) = "000000000000000000" else
       "00000000000000011000000000000000" when b(31 downto 15) = "00000000000000000" else
       "00000000000000001100000000000000" when b(31 downto 16) = "0000000000000000" else
       "00000000000000000110000000000000" when b(31 downto 17) = "000000000000000" else
       "00000000000000000011000000000000" when b(31 downto 18) = "00000000000000" else
       "00000000000000000001100000000000" when b(31 downto 19) = "0000000000000" else
       "00000000000000000000110000000000" when b(31 downto 20) = "000000000000" else
       "00000000000000000000011000000000" when b(31 downto 21) = "00000000000" else
       "00000000000000000000001100000000" when b(31 downto 22) = "0000000000" else
       "00000000000000000000000110000000" when b(31 downto 23) = "000000000" else
       "00000000000000000000000011000000" when b(31 downto 24) = "00000000" else
       "00000000000000000000000001100000" when b(31 downto 25) = "0000000" else
       "00000000000000000000000000110000" when b(31 downto 26) = "000000" else
       "00000000000000000000000000011000" when b(31 downto 27) = "00000" else
       "00000000000000000000000000001100" when b(31 downto 28) = "0000" else
       "00000000000000000000000000000110" when b(31 downto 29) = "000" else
       "00000000000000000000000000000011" when b(31 downto 30) = "00" else
       "00000000000000000000000000000001" when b(31)           = '0' else
       "00000000000000000000000000000000";
 
end architecture default;

